// IEEE 802.3-2022 82.2.8
// 40GBASE-R lane synchronization and reorderer
// delays blocks on each lane to align markers
// and reorders lanes based on marker data

module lane_deskew (
  input  logic clk,
  input  logic reset
);

endmodule : lane_deskew
