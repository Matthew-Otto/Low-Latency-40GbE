module eth_40gb (
  input logic
);

endmodule : eth_40gb
